// Module initialization
module inverter(
  input   a,      // input declaration
  output  y       // output declaration
);
  assign y = ~a;  // Assigning output value
endmodule
