module hello ();
	initial
		$display("hello I am Icarus");

endmodule
